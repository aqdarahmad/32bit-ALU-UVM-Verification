
// alu_subscriber.sv 
// Basic subscriber with simple coverage

class alu_subscriber extends uvm_subscriber #(alu_sequence_item);
  

  // Factory Registration

  `uvm_component_utils(alu_subscriber)
  

  // Transaction Handle

  alu_sequence_item sub;
  

  // Coverage Group
 
  covergroup aluCoverage;
    A: coverpoint sub.A;
    B: coverpoint sub.B;
    Opcode: coverpoint sub.Opcode;
    Result: coverpoint sub.Result;
    Error: coverpoint sub.Error;
  endgroup
  

  // Constructor

  function new(string name, uvm_component parent);
    super.new(name, parent);
    aluCoverage = new();
    sub = new();
  endfunction : new
  
 
  // Write Function

  function void write(alu_sequence_item t);
    sub.A = t.A;
    sub.B = t.B;
    sub.Opcode = t.Opcode;
    sub.Result = t.Result;  
    sub.Error = t.Error;
    aluCoverage.sample();
  endfunction : write
  

  // Report Phase

  function void report_phase(uvm_phase phase);
    super.report_phase(phase);
    `uvm_info(get_type_name(), 
              $sformatf("Coverage: %0.2f%%", aluCoverage.get_coverage()), 
              UVM_LOW)
  endfunction : report_phase
  
endclass : alu_subscriber